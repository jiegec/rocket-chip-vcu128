../../build/vcu128.RocketConfig.sv