../build/vcu128.SimConfig.sv